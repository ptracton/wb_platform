//                              -*- Mode: Verilog -*-
// Filename        : dsp_equations_sm.v
// Description     : DSP Equations State Machine
// Author          : Phil Tracton
// Created On      : Tue Apr 23 17:03:42 2019
// Last Modified By: Phil Tracton
// Last Modified On: Tue Apr 23 17:03:42 2019
// Update Count    : 0
// Status          : Unknown, Use with caution!
module dsp_equations_sm (/*AUTOARG*/
   // Inputs
   wb_clk, wb_rst
   ) ;
   input wb_clk;
   input wb_rst;

endmodule // dsp_equations_sm
